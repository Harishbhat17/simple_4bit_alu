module risc_5 #(parameter n=4)(input clk,

);